`define BR_BUS_LEN 34
`define IF_to_ID_LEN 64
`define ID_to_EXE_LEN 163
`define RF_BUS_LEN 38
`define EXE_to_MEM_LEN 109
`define MEM_to_WB_LEN 103
`define EXE_RF_LEN 38
`define MEM_RF_LEN 38
`define WB_RF_LEN  38
`define DEST_LEN 5

`define ST_W 7
`define ST_B 6
`define ST_H 5
`define LD_W 4
`define LD_B 3
`define LD_H 2
`define LD_BU 1
`define LD_HU 0

`define CSR_CRMD        3'h0
`define CSR_PRMD        3'h1
`define CSR_EUEN        3'h2
`define CSR_ECFG        3'h4
`define CSR_ESTAT       3'h5
`define CSR_ERA         3'h6
`define CSR_BADV        3'h7
`define CSR_EENTRY      3'hc
`define CSR_TLBIDX      3'h10
`define CSR_TLBEHI      3'h11
`define CSR_TLBELO0     3'h12
`define CSR_TLBELO1     3'h13
`define CSR_ASID        3'h18
`define CSR_PGDL        3'h19
`define CSR_PGDH        3'h1a
`define CSR_PGD         3'h1b
`define CSR_CPUID       3'h20
`define CSR_SAVE0       3'h30
`define CSR_SAVE1       3'h31
`define CSR_SAVE2       3'h32
`define CSR_SAVE3       3'h33
`define CSR_TID         3'h40
`define CSR_TCFG        3'h41
`define CSR_TVAL        3'h42
`define CSR_TICLR       3'h44
`define CSR_LLBCTL      3'h60
`define CSR_TLBRENTRY   3'h88
`define CSR_CTAG        3'h98
`define CSR_DMW0        3'h180
`define CSR_DMW1        3'h181

`define ECODE_INT   2'h0
`define ECODE_PIL   2'h1
`define ECODE_PIS   2'h2
`define ECODE_PIF   2'h3
`define ECODE_PME   2'h4
`define ECODE_PPI   2'h7
`define ECODE_ADE   2'h8
`define ECODE_ALE   2'h9
`define ECODE_SYS   2'hb
`define ECODE_BRK   2'hc
`define ECODE_INE   2'hd
`define ECODE_IPE   2'he
`define ECODE_FPD   2'hf
`define ECODE_FPE   2'h12
`define ECODE_TLBR  2'h3f

`define ESUBCODE_ADEF 1'b0
`define ESUBCODE_ADEM 1'b1